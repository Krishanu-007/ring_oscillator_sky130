** sch_path: /home/krishanu/Desktop/ring_oscillator_sky130/Xschem/Ring_Osc_3.sch
**.subckt Ring_Osc_3 Out
*.opin Out
x1 net4 Out net1 net3 inv
x2 net4 net1 net2 net3 inv
x3 net4 net2 Out net3 inv
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/krishanu/Desktop/ring_oscillator_sky130/Xschem/inv.sym
** sch_path: /home/krishanu/Desktop/ring_oscillator_sky130/Xschem/inv.sch
.subckt inv Vdd Vin Vout Vss
*.ipin Vin
*.ipin Vss
*.ipin Vdd
*.opin Vout
XM1 Vout Vin Vss GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vin Vdd VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
