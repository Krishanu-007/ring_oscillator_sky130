** RO_3_TEST flat netlist
*.OPIN OUT
*--------BEGIN_X1->RING_OSC_3
*.OPIN OUT
*.IPIN VSS
*.IPIN VDD
*.IPIN C1_-VE
*.IPIN C1_+VE
*.IPIN C2_-VE
*.IPIN C2_+VE
*.IPIN C3_+VE
*.IPIN C3_-VE
*--------BEGIN_X1_X1->INV
*.IPIN VIN
*.IPIN VSS
*.IPIN VDD
*.OPIN VOUT
*--------BEGIN_X1_X1_XM1->SKY130_FD_PR__NFET_01V8
XM1_X1_X1 NET1 OUT GND GND  SKY130_FD_PR__NFET_01V8 L=0.15 W=1 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29' PD='2*INT((NF+1)/2)*(W/NF+0.29)'
+ PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0 SD=0 MULT=1 M=1
*--------END___X1_X1_XM1->SKY130_FD_PR__NFET_01V8
*--------BEGIN_X1_X1_XM2->SKY130_FD_PR__PFET_01V8
XM2_X1_X1 NET1 OUT VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.15 W=2.5 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29' PD='2*INT((NF+1)/2)*(W/NF+0.29)'
+ PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0 SD=0 MULT=1 M=1
*--------END___X1_X1_XM2->SKY130_FD_PR__PFET_01V8
*--------END___X1_X1->INV
*--------BEGIN_X1_X2->INV
*.IPIN VIN
*.IPIN VSS
*.IPIN VDD
*.OPIN VOUT
*--------BEGIN_X1_X2_XM1->SKY130_FD_PR__NFET_01V8
XM1_X1_X2 NET6 NET1 GND GND  SKY130_FD_PR__NFET_01V8 L=0.15 W=1 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29' PD='2*INT((NF+1)/2)*(W/NF+0.29)'
+ PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0 SD=0 MULT=1 M=1
*--------END___X1_X2_XM1->SKY130_FD_PR__NFET_01V8
*--------BEGIN_X1_X2_XM2->SKY130_FD_PR__PFET_01V8
XM2_X1_X2 NET6 NET1 VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.15 W=2.5 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29' PD='2*INT((NF+1)/2)*(W/NF+0.29)'
+ PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0 SD=0 MULT=1 M=1
*--------END___X1_X2_XM2->SKY130_FD_PR__PFET_01V8
*--------END___X1_X2->INV
*--------BEGIN_X1_X3->INV
*.IPIN VIN
*.IPIN VSS
*.IPIN VDD
*.OPIN VOUT
*--------BEGIN_X1_X3_XM1->SKY130_FD_PR__NFET_01V8
XM1_X1_X3 OUT NET6 GND GND  SKY130_FD_PR__NFET_01V8 L=0.15 W=1 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29' PD='2*INT((NF+1)/2)*(W/NF+0.29)'
+ PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0 SD=0 MULT=1 M=1
*--------END___X1_X3_XM1->SKY130_FD_PR__NFET_01V8
*--------BEGIN_X1_X3_XM2->SKY130_FD_PR__PFET_01V8
XM2_X1_X3 OUT NET6 VDD VDD  SKY130_FD_PR__PFET_01V8 L=0.15 W=2.5 NF=1 AD='INT((NF+1)/2)*W/NF*0.29' AS='INT((NF+2)/2)*W/NF*0.29' PD='2*INT((NF+1)/2)*(W/NF+0.29)'
+ PS='2*INT((NF+2)/2)*(W/NF+0.29)' NRD='0.29/W' NRS='0.29/W' SA=0 SB=0 SD=0 MULT=1 M=1
*--------END___X1_X3_XM2->SKY130_FD_PR__PFET_01V8
*--------END___X1_X3->INV
*--------END___X1->RING_OSC_3
C1 NET1 NET2 10F M=1
C2 NET7 NET3 10F M=1
C3 NET5 NET4 10F M=1
C4 NET5 NET4 10F M=1
VDD VDD GND 1.8
**** BEGIN USER ARCHITECTURE CODE

.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt
.IC V(OUT)=0.01
.TRAN 100PS 10NS
.OPTIONS RELTOL=1E-4 ABSTOL=1E-12 VNTOL=1E-6
.SAVECURRENT
.SAVE ALL
.END

**** END USER ARCHITECTURE CODE
.end
